// ------------------------ Disclaimer -----------------------
// No warranty of correctness, synthesizability or 
// functionality of this code is given.
// Use this code under your own risk.
// When using this code, copy this disclaimer at the top of 
// Your file
//
// (c) Luca Hanel 2020
//
// ------------------------------------------------------------
//
// Module name: apb_bar
// 
// Functionality: Interconnect for APB bus
//
// Tests: 
//
// ------------------------------------------------------------

module apb_bar#(
  parameter APB_DATA_WIDTH = 32,
  parameter APB_ADDR_WIDTH = 32
)(

);

endmodule